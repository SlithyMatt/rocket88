// Rocket88 - A New 8-Bit Architecture
// Module: r88_alu
// Description: Arithmetic-Logic Unit
// See https://github.com/SlithyMatt/rocket88 for current code and documentation

module r88_alu(
 	input sysClock,
	inout [7:0] intD,
	input [7:0] regRight,
	input [7:0] regLeft,
	input [2:0] aluOp,
	input carryIn,
	output carryOut,
	input invOut,
	input decMode,
	input carryInEn,
	input rightSel
);


endmodule
